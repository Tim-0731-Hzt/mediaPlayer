--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   14:44:00 10/07/2020
-- Design Name:   
-- Module Name:   C:/Users/seanw/Local Documents/UNSW/COMP3601/COMP3601/VHDL/IR_Decoder_Testbench.vhd
-- Project Name:  IR_Decoder
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: IR_Decoder
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY IR_Decoder_Testbench IS
END IR_Decoder_Testbench;
 
ARCHITECTURE behavior OF IR_Decoder_Testbench IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT IR_Decoder
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         ir : IN  std_logic;
         data : OUT  std_logic_vector(11 downto 0);
         done : OUT  std_logic
        );
    END COMPONENT;
	
	COMPONENT Timer
    PORT(
         clk : IN  std_logic;
         en : IN  std_logic;
         reset : IN  std_logic;
         usec : INOUT  integer;
         msec : INOUT  integer
        );
    END COMPONENT;

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal ir : std_logic := '1';

 	--Outputs
   signal data : std_logic_vector(11 downto 0);
   signal done : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: IR_Decoder PORT MAP (
          clk => clk,
          reset => reset,
          ir => ir,
          data => data,
          done => done
        );
		

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
	  
      wait for clk_period*10;
		reset <= '1';
      ir <= '0';

      wait for 2700 us;
      -- insert stimulus here 
		ir <= '1';
		
	wait for 100 us;
	
		ir <= '0';
		
	wait for 600 us;
		ir <= '1';
      wait;
   end process;

END;
